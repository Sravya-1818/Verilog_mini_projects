module gray_code(y,a);
  output [3:0]y;
  input [3:0]a;
  assign y[3]=a[3];
  assign y[2]=a[3]^a[2];
  assign y[1]=a[2]^a[1];
  assign y[0]=a[1]^a[0];
endmodule
